module bikeTrailEdge(bikeLocation_middle, vga_address, bike_orient, trail_over_bike);
	input [18:0] bikeLocation_middle;
	input [18:0] vga_address;
	input [1:0] bike_orient;
	output trail_over_bike;
	
	
endmodule