/**
 * The processor takes in two inputs and returns two outputs
 *
 * Inputs
 * clock: this is the clock for your processor at 50 MHz
 * reset: we should be able to assert a reset to start your pc from 0 (sync or
 * async is fine)
 *
 * Outputs
 * dmem_data_in: this should connect to the wire that feeds in data to your dmem
 * dmem_address: this should be the address of data that you write data to
 *
 * Notes
 * You will need to figure out how to instantiate two memory elements, called
 * "syncram," in Quartus: one for imem and one for dmem. Each should take in a
 * 12-bit address and allow for storing a 32-bit value at each address. Each
 * should have a single clock.
 *
 * Each memory element should have a corresponding .mif file that initializes
 * the memory element to certain value on start up. These should be named
 * imem.mif and dmem.mif respectively.
 *
 * imem
 * Inputs:  12-bit address, 1-bit clock enable, and a clock
 * Outputs: 32-bit instruction
 *
 * dmem
 * Inputs:  12-bit address, 1-bit clock, 32-bit data, 1-bit write enable
 * Outputs: 32-bit data at the given address
 *
 */ 
module processor(masterSwitch, clock, reset, dmem_data_in, dmem_address, instructionFDout, pcout, pcFDout, pcDXout, pcXMout, j1enDXout, j2enDXout, ren_outDXout, ren_outXMout, ren_outMWout, menDXout, benDXout, exenDXout, OoutXMout, BoutXMout, aluopDXout, aluopfin, shamtDXout, rd_outDXout, ADXout, BDXout, selectDXout, selectXMout, dataMWout, OoutMWout, selectMWout, rd_outXMout, rd_outMWout, readADXout, readBDXout, readBXMout, dataW, readAD, readBD, stall, flush, benfinal, bikeblue, bikeblueOrient,reg27);
    input clock, reset, masterSwitch;

    output [31:0] dmem_data_in;
    output [11:0] dmem_address;
	 
	 assign dmem_data_in = datawritefinal;
	 assign dmem_address = OoutXMout[11:0]; 
	 
	 // Instantiate all outputs from D
	 wire j1enDin, j2enDin, ren_outDin, menDin, benDin, exenDin;
	 wire j1enDout, j2enDout, ren_outDout, menDout, benDout, exenDout;
	 dffe1 j1d_dff(.d(j1enDin),.q(j1enDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));  // J1D
	 dffe1 j2d_dff(.d(j2enDin),.q(j2enDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));  // J2D
	 dffe1 rend_dff(.d(ren_outDin),.q(ren_outDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Ren_out D
	 dffe1 mend_dff(.d(menDin),.q(menDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));   // MD
	 dffe1 bend_dff(.d(benDin),.q(benDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));   // BD
	 dffe1 exend_dff(.d(exenDin),.q(exenDout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // ED	
	 
	 // Instantiate all outputs from DX
	 output j1enDXout, j2enDXout, ren_outDXout, menDXout, benDXout, exenDXout;
	 dffe1 j1dx_dff(.d(j1enDout),.q(j1enDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));  // J1DX
	 dffe1 j2dx_dff(.d(j2enDout),.q(j2enDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));  // J2DX
	 dffe1 rendx_dff(.d(ren_outDout),.q(ren_outDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Ren_out DX
	 dffe1 mendx_dff(.d(menDout),.q(menDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));   // MDX
	 dffe1 bendx_dff(.d(benDout),.q(benDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));   // BDX
	 dffe1 exendx_dff(.d(exenDout),.q(exenDXout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // EDX
	 
	 // Need to be passed on to execute
	 output ren_outXMout;
	 wire ren_outXout;
	 dffe1 renx_dff(.d(ren_outDXout),.q(ren_outXout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
	 dffe1 renxm_dff(.d(ren_outXout),.q(ren_outXMout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Ren_out, XM	 
	 
	 // Need to be passed on to memory
	 wire ren_outMout;
	 output ren_outMWout;
	 dffe1 renm_dff(.d(ren_outXMout),.q(ren_outMout),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
	 dffe1 renmw_dff(.d(ren_outMout),.q(ren_outMWout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Ren_out, XM
	 
	 output [4:0] shamtDXout, aluopDXout, rd_outDXout;
	 wire [4:0] shamtDXin, aluopDXin, rd_outDXin, readADout, readBDout, readBXout;
	 wire [4:0] shamtDin, aluopDin, rd_outDin, rd_outXin, readADin, readBDin, shamtDout, aluopDout, rd_outDout, rd_outXout, rd_outMout, rd_outWout;
	 output [4:0] rd_outXMout, rd_outMWout, readADXout, readBDXout, readBXMout;
	 genvar h;
	 generate
		for(h=0;h<5;h=h+1) begin : Hloop
			dffe1 readAD_dff(.d(readADin[h]),.q(readADout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));  //Used for Bypasses in X
			dffe1 readADX_dff(.d(readADout[h]),.q(readADXout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); 
			
			dffe1 readBD_dff(.d(readBDin[h]),.q(readBDout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 readBDX_dff(.d(readBDout[h]),.q(readBDXout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 readBX_dff(.d(readBDXout[h]),.q(readBXout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 readBXM_dff(.d(readBXout[h]),.q(readBXMout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			
			dffe1 shamtd_dff(.d(shamtDin[h]),.q(shamtDout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 shamtdx_dff(.d(shamtDout[h]),.q(shamtDXout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			
			dffe1 aluop_dff(.d(aluopDin[h]),.q(aluopDout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));			
			dffe1 aluopdx_dff(.d(aluopDout[h]),.q(aluopDXout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			
			dffe1 rd_outD_dff(.d(rd_outDin[h]),.q(rd_outDout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 rd_outDX_dff(.d(rd_outDout[h]),.q(rd_outDXout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 rd_outX_dff(.d(rd_outXin[h]),.q(rd_outXout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 rd_outXM_dff(.d(rd_outXout[h]),.q(rd_outXMout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 rd_outM_dff(.d(rd_outXMout[h]),.q(rd_outMout[h]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 rd_outMW_dff(.d(rd_outXMout[h]),.q(rd_outMWout[h]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
		end
	 endgenerate	
	 
	 output [11:0] pcout, pcFDout, pcDXout, pcXMout;
	 wire [11:0] pcDout, pcXout, pcXin, pcXMin, pcin;
	 genvar i;
	 generate
		for(i=0;i<12;i=i+1) begin : PCloop
		   dffe1 pc_dff(.d(pcin[i]),.q(pcout[i]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // PC
			dffe1 pcfd_dff(.d(pcout[i]),.q(pcFDout[i]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // F/D
			dffe1 pcd_dff(.d(pcFDout[i]),.q(pcDout[i]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // D
			dffe1 pcdx_dff(.d(pcDout[i]),.q(pcDXout[i]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // D/X
			dffe1 pcx_dff(.d(pcDXout[i]),.q(pcXout[i]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // X
			dffe1 pcxm_dff(.d(pcXout[i]),.q(pcXMout[i]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // X/M
		end
	 endgenerate
	 
	 wire [16:0] immediateDXin, immediateDin, immediateDout;
	 wire [16:0] immediateDXout;
	 genvar k;
	 generate
		for(k=0;k<17;k=k+1) begin:Loop17
			dffe1 imm_dff(.d(immediateDin[k]),.q(immediateDout[k]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 immdx_dff(.d(immediateDout[k]),.q(immediateDXout[k]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
		end
	 endgenerate
	 
	 wire [26:0] targetDXin, targetDin, targetDout;
 	 wire [26:0] targetDXout;
	 genvar l;
	 generate
		for(l=0;l<27;l=l+1) begin: Loop27
			dffe1 targetd_dff(.d(targetDin[l]),.q(targetDout[l]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
			dffe1 targetdx_dff(.d(targetDout[l]),.q(targetDXout[l]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
		end
	 endgenerate
	 
	 output [31:0] instructionFDout, OoutXMout, BoutXMout, ADXout, BDXout, selectDXout, selectXMout, selectMWout, dataMWout, OoutMWout, dataW;
	 wire [31:0] instructionFDin, OoutXMin, BoutXMin;
	 wire [31:0] ADXin, BDXin, selectDXin, selectXMin, selectMWin, dataMWin, dataWBin;
	 wire [31:0] ADin, BDin, selectDin, selectXin, OoutXin, BoutXin, ADout, BDout, selectDout, selectXout, selectMout, OoutXout, BoutXout, OoutMout;
	 genvar j;
	 generate 
		for(j=0;j<32;j=j+1) begin: Loop32
			dffe1 inst_dff(.d(instructionFDin[j]),.q(instructionFDout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Instruction in latch F/D
	
			dffe1 select_Ddff(.d(selectDin[j]),.q(selectDout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch D
			
			dffe1 ADX_dff(.d(ADXin[j]),.q(ADXout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // A in latch D/X
			dffe1 BDX_dff(.d(BDXin[j]),.q(BDXout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // B in latch D/X
			dffe1 selectDX_dff(.d(selectDout[j]),.q(selectDXout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch D/X
			
			dffe1 selectX_dff(.d(selectDXout[j]),.q(selectXout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch X
			dffe1 OoutX_dff(.d(OoutXin[j]),.q(OoutXout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Oout in X latch
			dffe1 BoutX_dff(.d(BoutXin[j]),.q(BoutXout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Bout in X latch
			
			dffe1 selectxm_dff(.d(selectXout[j]),.q(selectXMout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch X/M
			dffe1 OoutXM_dff(.d(OoutXout[j]),.q(OoutXMout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Oout in XM latch
			dffe1 BoutXM_dff(.d(BoutXout[j]),.q(BoutXMout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Bout in XM latch
			
			dffe1 selectm_dff(.d(selectXMout[j]),.q(selectMout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch M
			dffe1 OoutM_dff(.d(OoutXMout[j]),.q(OoutMout[j]),.clk(~clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Oout in M latch
			
			dffe1 selectmw_dff(.d(selectMout[j]),.q(selectMWout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Select in latch M/W
			dffe1 OoutMW_dff(.d(OoutMout[j]),.q(OoutMWout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Oout in MW latch
			dffe1 dataMWout_dff(.d(dataMWin[j]),.q(dataMWout[j]),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1)); // Data out in MW latch
			end
	 endgenerate
	 
	 output stall;
	 
	 // Choose where the next PC is
	 wire firstin, firstout;
	 output flush;
	 dffe1 first_dffe(.d(firstin),.q(firstout),.clk(clock),.ena(1'b1),.clrn(~reset),.prn(1'b1));
	 pc mypc(.next(pcin),.current(pcout), .stall(stall), .prev(pcFDout), .reset(reset), .jump1en(j1enDXout), .jump2en(j2enDXout), .ben(benfinal),.jumprt(ADXout[11:0]), .jumpt(targetDXout[11:0]),.N(immediateDXout), .firstin(firstout), .firstout(firstin),.flush(flush));
	 
	 // Fetch
	 F myF(.clock(clock),.pcin(pcin),.instruction(instructionFDin));
	 
	 // Stall Logic
	 output[4:0] readAD, readBD;
	 stall mystall(stall, selectDXout[8], rd_outDXout, instructionFDout, j1enDin, j2enDin, ren_outDin, menDin, benDin, exenDin, aluopDin, shamtDin, rd_outDin, readAD, readBD, immediateDin, targetDin, selectDin, flush);	 
	 assign readADin = readAD;
	 assign readBDin = readBD;
	 
	 // Decode
	 output [31:0] bikeblue, bikeblueOrient;
	 output reg27;
	 D myD(ADXin, BDXin, readAD, readBD, clock, reset, ren_outMWout, rd_outMWout, dataW, bikeblue, bikeblueOrient, masterSwitch, reg27);
	 
	 
	 // eXecute
	 output [4:0] aluopfin;
	 output benfinal;
	 X myX(menDXout, benDXout, exenDXout, aluopDXout, ADXout, BDXout, readADXout, readBDXout, rd_outDXout, rd_outXin, ren_outXMout, rd_outXMout, OoutXMout, ren_outMWout, rd_outMWout, dataW, selectDXout, immediateDXout, targetDXout, shamtDXout, aluopfin, OoutXin, BoutXin, reset, pcDXout, benfinal);	 
	 
	 // Memory, BoutXMout is rd data, OoutXMout is rs+N address (or should be)
	 wire [31:0] datawritefinal;
	 M myM(.swen(selectXMout[7]),.clock(clock), .data_write(BoutXMout), .data_where(OoutXMout), .data_mem(dataMWin), .readXM(readBXMout), .renWB(ren_outMWout), .readWB(rd_outMWout), .dataWB(dataW), .data_writefinal(datawritefinal));
	 
	 // WriteBack
	 W myW(dataMWout,OoutMWout,selectMWout[8],dataW);
	 
endmodule

